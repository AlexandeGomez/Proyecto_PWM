module controlDireccion(
output in1, in2
);

assign in1 = 1'b1;
assign in2 = 1'b0;

endmodule
